/* 
  This is my LEF!
*/
